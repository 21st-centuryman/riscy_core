`timescale 10ns/1ns

module TB();
  // ADD INPUTS
  
  ALU DUT(OP,A,B, ONZ, Result); // EDIT THIS

  initial begin
   // Add
  end
endmodule
